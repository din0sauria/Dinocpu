`timescale 1ns / 1ps
//顶层模块负责连接系统核心组件（CPU、存储、时钟、IO），通过内部信号（wire）传递控制与数据
//最终实现「指令执行-数据存储-状态显示」的完整流程，并支持通过开关（sw_i）进行调试控制。
module PLCPUSOC_Top(
        input   clk,
        input   rstn,
        input  [15:0] sw_i, // output to switch
        output [7:0] disp_seg_o, disp_an_o // output to seg7
   );
  
   wire Clk_CPU;        // CPU clock
   wire [31:0]  instr;  // instruction
   wire [31:0]  pc;     // PC
   wire memwrite;       // memory write
   wire memread;        // memory read        new add
   wire [31:0]  dm_din, dm_dout; // data 
   
   wire rst;
   assign rst = ~rstn;

   wire [31:0] seg7_data; 
   wire [6:0]  ram_addr;
   wire ram_we;
   wire seg7_we;
   
   wire [31:0]  cpu_data_out;       // data from CPU
   wire [31:0]  cpu_data_addr;
   wire [31:0]  ram_data_out;
   wire [31:0]  cpu_data_in;
   wire [31:0]  cpuseg7_data;
   wire [31:0]  reg_data;
   
  // 时钟管理
   clk_div U_CLKDIV( 
         .clk(clk),       // board clock
         .rst(rst),       // reset 
         .SW15(sw_i[15]), // sw15
         .Clk_CPU(Clk_CPU)// cpu clock
         );
         
  // instantiation of single-cycle cpu       
   PLCPU U_PLCPU(
         .clk(Clk_CPU),             // cpu clock
         .reset(rst),               // reset
         .inst_in(instr),           // instruction
         .Data_in(cpu_data_in),     // data from meory/IO to cpu  
         .mem_w(memwrite),          // memory/IO(seg7) write signal
         .mem_r(memread),           // memory/IO(seg7) read signal   new add signal
         .PC_out(pc),               // PC
         .Addr_out(cpu_data_addr),  // address from cpu to memory/IO(seg7)
         .Data_out(cpu_data_out),   // data from cpu to memory/IO
         .reg_sel(sw_i[4:0]),       // register selection
         .reg_data(reg_data)        // register data
         );

  // instantiation of intruction memory (used for FPGA), imem is generated by IP core
  //存储系统
  //指令存储器
   imem  U_IM(
         .a(pc[8:2]), .spo(instr)
         );

  //数据存储器
   dm    U_DM(
         .clk(Clk_CPU),   // cpu clock
         .DMWr(ram_we),   // ram write
         .DMRe(memread),                // new add
         .addr({23'b0, ram_addr, 2'b00}), // ram address
         .din(dm_din),    // data to ram
         .dout(dm_dout)   // data from ram
         );

  // 总线与 IO 管理
   MIO_BUS  U_MIO (
         .sw_i(sw_i),                   // switch
         .mem_w(memwrite),              // memory/IO(seg7) write signal
         .cpu_data_out(cpu_data_out),   // data from cpu to memory/IO 
         .cpu_data_addr(cpu_data_addr), // address from cpu to memory/IO(seg7)
         .ram_data_out(dm_dout),        // data from ram 
         .cpu_data_in(cpu_data_in),     // data from memory/IO to cpu
         .ram_data_in(dm_din),          // data to ram
         .ram_addr(ram_addr),           // ram address
         .cpuseg7_data(cpuseg7_data),   // data from cpu to seg7
         .ram_we(ram_we),               // memory write signal
         .seg7_we(seg7_we)              // seg7 write signal
   );
   
  // 状态显示（Multi_CH32 + seg7x16）
  //Multi_CH32（多路选择器）：通过开关 sw_i[5:0] 选择 8 个调试通道（如 PC、指令、地址、内存数据等），输出待显示的 seg7_data。
   Multi_CH32 U_Multi (
          .clk(clk),                        // board clk
          .rst(rst),                        // reset
          .EN(seg7_we),                     // seg7 write enable
          .ctrl(sw_i[5:0]),                 // SW[5:0]
          .Data0(cpuseg7_data),             // channel 0 (data from cpu to seg7)
           //disp_cpudata
          .data1({2'b0,pc[31:2]}),          // test channel 1--instruction no.
          .data2(pc),                       // test channel 2--PC
          .data3(instr),                    // test channel 3--instruction
          .data4(cpu_data_addr),            // test channel 4--address from cpu to memory/IO(seg7)
          .data5(cpu_data_out),             // test channel 5--data from cpu to memory/IO
          .data6(dm_dout),                  // test channel 6--data from ram
          .data7({23'b0, ram_addr, 2'b00}), // test channel 7--ram address
          .reg_data(reg_data),              // selected register data
          .seg7_data(seg7_data)             // data to seg7 display
          );
            
  // seg7x16（数码管驱动）：将 seg7_data 转换为实际硬件的段选（disp_seg_o）和位选（disp_an_o）信号，驱动 16 位数码管显示系统状态（支持调试观察）。       
   seg7x16 U_7SEG(
         .clk(clk),           // board clock
         .rst(rst),           // reset
         .cs(1'b1),           // selection (always 1)
         .i_data(seg7_data),  // data to seg7 display
         .o_seg(disp_seg_o),  // to board disp_seg_o
         .o_sel(disp_an_o)    // to board disp_an_o
         );

endmodule
